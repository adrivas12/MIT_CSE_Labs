module q4(G, L, E, x,y);
	input [4:0] a, b;
	output G, L, E;
	E = (~(a[4]^b[4]))&(~(a[3]^b[3]))&(~(a[2]^b[2]))&(~(a[1]&b[1]))&(~(a[0]^b[0]));
	G = (a[4]&~b[4])|((~(a[4]^b[4]))&(a[3]&b[3]))|(~(a[4]^b[4])&(~(a[3]^b[3]))&(a[2]&~b[2])) | ((~(a[4]^b[4]))&(~(a[3]^b[3]))&(~(a[2]^b[2]))&(a[1]&~b[1]))|(~(a[4]^b[4])&(~(a[3]^b[3]))&(~(a[2]^b[2]))&(~(a[1]&b[1]))&(a[0]&~b[0]))

	L=(~a[4]&b[4])|((~(a[4]^b[4]))&(a[3]&b[3]))|(~(a[4]^b[4])&(~(a[3]^b[3]))&(a[2]&~b[2]))|(~(a[4]^b[4])&(~(a[3]^b[3]))&(~(a[2]^b[2]))&(a[1]&~b[1]))|((a[4]&~b[4])&(~(a[3]^b[3]))&(~(a[2]^b[2]))&(~(a[1]&b[1]))&(a[0]&~b[0]))