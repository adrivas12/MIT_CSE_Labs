`timescale 1ns/1ns
`include "q5.v"

module q5_tb();
reg [0:15]W;
wire [0:3]Y;
wire Z;
q5 q5(W, Z, Y);
initial 
begin

	$dumpfile("q5_tb.vcd");
	$dumpvars(0, q5_tb);

	W=16'b 1000000000000000; #10;
	W=16'b 0100000000000000; #10;
	W=16'b 0010000000000000; #10;
	W=16'b 0001000000000000; #10;
	W=16'b 0000100000000000; #10;
	W=16'b 0000010000000000; #10;
	W=16'b 0000001000000000; #10;
	W=16'b 0000000100000000; #10;
	W=16'b 0000000010000000; #10;
	W=16'b 0000000001000000; #10;
	W=16'b 0000000000100000; #10;
	W=16'b 0000000000010000; #10;
	W=16'b 0000000000001000; #10;
	W=16'b 0000000000000100; #10;
	W=16'b 0000000000000010; #10;
	W=16'b 0000000000000001; #10;


	$display("Test Completed");

end 
endmodule