`timescale 1ns/1ns
`include "q3.v"

module q3_tb();
reg [15:0]w;
reg [3:0]s;
wire f;

q3 q3(w, s, f);
initial 
begin
	$dumpfile("q3_tb.vcd");
	$dumpvars(0,q3_tb);

	w=16'b0001110001110001; s=4'b0000;
	#10;
	w=16'b0001110001110001; s=4'b0001;
	#10;
	w=16'b0001110001110001; s=4'b0010;
	#10;
	w=16'b0001110001110001; s=4'b0011;
	#10;
	w=16'b0001110001110001; s=4'b0100;
	#10;
	w=16'b0001110001110001; s=4'b0101;
	#10;
	w=16'b0001110001110001; s=4'b0110;
	#10;
	w=16'b0001110001110001; s=4'b0111;
	#10;
	w=16'b0001110001110001; s=4'b1000;
	#10;
	w=16'b0001110001110001; s=4'b1001;
	#10;
	w=16'b0001110001110001; s=4'b1010;
	#10;
	w=16'b0001110001110001; s=4'b1011;
	#10;
	w=16'b0001110001110001; s=4'b1100;
	#10;
	w=16'b0001110001110001; s=4'b1101;
	#10;
	w=16'b0001110001110001; s=4'b1110;
	#10;
	w=16'b0001110001110001; s=4'b1111;
	#10;

	$display("test complete");
end
endmodule